`ifndef __PIPES_SV
`define __PIPES_SV

package pipes;
    import common::*;
    
/* Define instruction decoding rules here */

// parameter F6_R_TYPE = 6'bxxxxxxx;

/* Define pipeline structures here */


endpackage

`endif
